`ifndef STB_DEC__SV
`define STB_DEC__SV

package stb_dec;
    
    parameter ON = 1;
    parameter OFF = 0;
    
endpackage
`endif
